��<N      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.2�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�auto�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�objawy��wiek��choroby_wsp��wzrost��leki�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh$hNhJ�
hG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��h2�f8�����R�(KhINNNJ����J����K t�b�C              �?�t�bhMh&�scalar���hHC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hK�
node_count�K�nodes�h(h+K ��h-��R�(KK��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hyhHK ��hzhHK��h{hHK��h|hYK��h}hYK ��h~hHK(��hhYK0��uK8KKt�b�B                            �<@�D����?             E@������������������������       �                     @                            @����X�?            �A@                          �E@      �?             8@                         ��e@���Q��?             @������������������������       �                     �?                          �@@      �?             @������������������������       �                     �?	       
                   �g@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @                          �Q@�}�+r��?             3@������������������������       �        
             .@                           S@      �?             @������������������������       �                     �?������������������������       �                     @                           @���|���?             &@                         ��g@      �?             @������������������������       �                     @������������������������       �                     �?                          �P@؇���X�?             @������������������������       �                     @������������������������       �                     �?�t�b�values�h(h+K ��h-��R�(KKKK��hY�Bp        9@      1@              @      9@      $@      5@      @      @       @              �?      @      �?      �?               @      �?      �?              �?      �?      2@      �?      .@              @      �?              �?      @              @      @      @      �?      @                      �?      �?      @              @      �?        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ/��hG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�BH         
                    �?և���X�?             E@       	                  y�E@և���X�?             <@                          Pd@�����H�?             2@������������������������       �                     �?                          �g@�IєX�?             1@������������������������       �                     (@                           @z�G�z�?             @������������������������       �                     @������������������������       �      �?              @������������������������       �                     $@                           �?؇���X�?	             ,@������������������������       �                     �?                          �C@$�q-�?             *@������������������������       �                     �?������������������������       �                     (@�t�bh�h(h+K ��h-��R�(KKKK��hY�C�      8@      2@      (@      0@       @      0@      �?              �?      0@              (@      �?      @              @      �?      �?      $@              (@       @              �?      (@      �?              �?      (@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJu�7hG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�Bx                            �E@և���X�?             E@       	                    @�r����?	             .@                            @$�q-�?             *@                          �5@z�G�z�?             @������������������������       �                     @                          �B@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @
                          �@@      �?              @������������������������       �                     �?������������������������       �                     �?                            @�+$�jP�?             ;@                           �?�����H�?
             2@������������������������       �                     "@                         y�H@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @                         �%g@�q�q�?             "@������������������������       �                     @                           �?      �?             @                            @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KKKK��hY�B�        8@      2@       @      *@      �?      (@      �?      @              @      �?      �?      �?                      �?               @      �?      �?              �?      �?              6@      @      0@       @      "@              @       @               @      @              @      @      @              @      @      @      �?      @                      �?               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��!XhG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�B�                              �?�G��l��?             E@                          �g@d}h���?	             ,@������������������������       �                     &@������������������������       �                     @                           0@��>4և�?             <@������������������������       �                      @                          `h@$��m��?             :@       	                   �:@�\��N��?             3@������������������������       �                      @
                           �?��.k���?             1@������������������������       �                     @                           @�	j*D�?	             *@������������������������       �                      @                          �P@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKKK��hY�B        6@      4@      &@      @      &@                      @      &@      1@       @              "@      1@      "@      $@               @      "@       @              @      "@      @       @              �?      @              @      �?                      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJC�NhG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�Bx                             @�q�q�?             E@       	                   @C@"pc�
�?             6@                            @���Q��?             @                           �?      �?             @                          `d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?
                           @�IєX�?             1@������������������������       �                     *@                          pf@      �?             @������������������������       �                     @������������������������       �                     �?                          �g@      �?             4@                          �@@      �?             (@������������������������       �                     �?                            @"pc�
�?             &@������������������������       �                     "@������������������������       �                      @                          �<@      �?              @������������������������       �                     @                          �g@z�G�z�?             @������������������������       �                      @������������������������       ��q�q�?             @�t�bh�h(h+K ��h-��R�(KKKK��hY�B�        <@      ,@      2@      @       @      @       @       @      �?       @      �?                       @      �?                      �?      0@      �?      *@              @      �?      @                      �?      $@      $@      "@      @              �?      "@       @      "@                       @      �?      @              @      �?      @               @      �?       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�R�[hG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�B(         
                  y�E@�ՙ/�?             E@                          Pd@�t����?             1@������������������������       �                     @                          �@@$�q-�?
             *@������������������������       �                      @       	                     @z�G�z�?             @                          �f@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �?�J�4�?             9@������������������������       �                     &@                          Ph@����X�?
             ,@                          @N@r�q��?	             (@                            @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KKKK��hY�B0        :@      0@      @      (@      @              �?      (@               @      �?      @      �?      �?              �?      �?                      @      5@      @      &@              $@      @      $@       @      @       @      @                       @      @                       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�v}hG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�B�                            �@@��6���?             E@                           0@$�q-�?             *@                         �ee@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@                           N@>���Rp�?             =@                            @��Q��?             4@	       
                   �d@d}h���?	             ,@������������������������       �                     �?                         y�H@8�Z$���?             *@                           @����X�?             @������������������������       �                     @                         y
F@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @                          �H@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@�t�bh�h(h+K ��h-��R�(KKKK��hY�BP        7@      3@      �?      (@      �?      �?      �?                      �?              &@      6@      @      *@      @      &@      @              �?      &@       @      @       @      @               @       @       @                       @      @               @      @       @                      @      "@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJg}�XhG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�B�         
                   �@@և���X�?             E@       	                     @�<ݚ�?             "@                           �?�q�q�?             @                          pd@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         �5g@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                           �?�q�q�?            �@@������������������������       �                     $@                           @
;&����?             7@                           �?X�Cc�?             ,@������������������������       �                      @                         y
N@�q�q�?             (@                          �E@�z�G��?             $@                            @      �?              @                           @����X�?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                          �N@�q�q�?             "@������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKKK��hY�B�        8@      2@       @      @       @      @      �?       @      �?                       @      �?       @      �?                       @              @      6@      &@      $@              (@      &@      "@      @       @              @      @      @      @      @      @      @       @      �?              @       @              �?       @                       @      @      @              @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ	�tlhG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�B�                             @�G��l��?             E@       	                  �%g@      �?             4@                            �?@4և���?	             ,@������������������������       �                     @                          �E@      �?              @                          �d@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @
                          0h@�q�q�?             @                            @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                         y�H@�X����?             6@                          �@@�t����?
             1@������������������������       �                      @                           @�<ݚ�?             "@                            @����X�?             @                          �g@���Q��?             @������������������������       �                     �?                         y�C@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKKK��hY�B�        6@      4@      .@      @      *@      �?      @              @      �?      @      �?      @                      �?      @               @      @      �?      @      �?                      @      �?              @      .@       @      .@               @       @      @       @      @       @      @      �?              �?      @      �?       @              �?               @               @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�ޡhG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�B(                           y�E@�G��l��?             E@       	                    @z�G�z�?             4@                          `d@      �?	             0@������������������������       �                     �?                          �;@��S�ۿ?             .@������������������������       �                     @                           �?      �?              @������������������������       �                     �?������������������������       �                     @
                          �g@      �?             @������������������������       �                      @������������������������       �                      @                          @N@"pc�
�?             6@                           �?�	j*D�?             *@������������������������       �                      @                          0f@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@�t�bh�h(h+K ��h-��R�(KKKK��hY�B0        6@      4@      @      0@       @      ,@      �?              �?      ,@              @      �?      @      �?                      @       @       @               @       @              2@      @      "@      @       @              �?      @      �?                      @      "@        �t�bubhhubehhub.